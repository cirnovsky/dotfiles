Vim�UnDo� �2~K���ȡ����Ɔ�=��b��S���      	                             h���    _�                             ����                                                                                                                                                                                                                                                                                                                                                             h���     �                   5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             h�ك     �                >module theormo(input [7:0] Tset, [7:0] Tact, output Hon, Con);    �                �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             h�ن     �                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�ُ     �                >module theormo(input [7:0] Tset, [7:0] Tact, output Hon, Con);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�ْ     �                Cmodule theormo #() (input [7:0] Tset, [7:0] Tact, output Hon, Con);5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             h�ٙ     �                Rmodule theormo #(parameter LEN=8) (input [7:0] Tset, [7:0] Tact, output Hon, Con);5�_�                       :    ����                                                                                                                                                                                                                                                                                                                                                             h�ٛ     �                Vmodule theormo #(parameter LEN=8) (input [LEN-1:0] Tset, [7:0] Tact, output Hon, Con);5�_�      	                 >    ����                                                                                                                                                                                                                                                                                                                                                             h�ٞ    �                Ymodule theormo #(parameter LEN=8) (input [LEN-1:0] Tset, [LEN-:0] Tact, output Hon, Con);5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                v       h�ٱ     �                Zmodule theormo #(parameter LEN=8) (input [LEN-1:0] Tset, [LEN-1:0] Tact, output Hon, Con);5�_�   	              
      ,    ����                                                                                                                                                                                                                                                                                                                               ,          .       v       h�ٴ     �                \module theormo #(parameter width=8) (input [LEN-1:0] Tset, [LEN-1:0] Tact, output Hon, Con);5�_�   
                    >    ����                                                                                                                                                                                                                                                                                                                               >          @       v   0    h�ٴ    �                ^module theormo #(parameter width=8) (input [width-1:0] Tset, [LEN-1:0] Tact, output Hon, Con);5�_�                           ����                                                                                                                                                                                                                                                                                                                               >          @       v   0    h���     �               	5�_�                           ����                                                                                                                                                                                                                                                                                                                               >          @       v   0    h���     �                `module theormo #(parameter width=8) (input [width-1:0] Tset, [width-1:0] Tact, output Hon, Con);    �                �             5�_�                           ����                                                                                                                                                                                                                                                                                                                               >          @       v   0    h���     �               	assign Hon = 5�_�                           ����                                                                                                                                                                                                                                                                                                                               >          @       v   0    h���     �                  �               5�_�                            ����                                                                                                                                                                                                                                                                                                                               >          @       v   0    h���    �               module jdoodle;    �                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        h��a     �                �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h��x     �                `module theormo #(parameter width=8) (input [width-1:0] Tset, [width-1:0] Tact, output Hon, Con);5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h��}     �                bmodule thermormo #(parameter width=8) (input [width-1:0] Tset, [width-1:0] Tact, output Hon, Con);5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h��}     �                amodule thermoro #(parameter width=8) (input [width-1:0] Tset, [width-1:0] Tact, output Hon, Con);5�_�                          ����                                                                                                                                                                                                                                                                                                                                         
       v       h�ڃ    �                `module thermor #(parameter width=8) (input [width-1:0] Tset, [width-1:0] Tact, output Hon, Con);5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h�ڄ     �   
            	thermo5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h�ڽ     �               	�             5�_�                            ����                                                                                                                                                                                                                                                                                                                                         
       v       h���     �               #1;5�_�                            ����                                                                                                                                                                                                                                                                                                                                         
       v       h���    �               #1;5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h���     �               		�             5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h���    �               	�             5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h���     �               	�             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V   
    h���    �               	Tset = 50;   	$display("Tset=%d", Tset);   	$display(" Tact | Hon Con");   	$display("----------------");       0	for (integer i = 40; i <= 60; i = i + 2) begin;   		Tact = i;   		#1;   .		$display(" %2d  | %b   %b", Tact, Hon, Con);   	end   		$finish;5�_�                           ����                                                                                                                                                                                                                                                                                                                                         
       v       h�ځ     �                _module thermor#(parameter width=8) (input [width-1:0] Tset, [width-1:0] Tact, output Hon, Con);5��